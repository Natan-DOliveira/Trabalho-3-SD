module tb_fila;

endmodule