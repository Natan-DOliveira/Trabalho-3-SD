module tb_fila;